`timescale 1ns / 1ps
module instance_module();
endmodule


module test_source();
    instance_module u_inst();
endmodule
